`timescale 1ns/1ns;

module TOP;



endmodule
